`timescale 1ns/1ns
module DataPath(
	clk,
	rst, 
	start_par,
    	start_rot, 
    	start_per,  
    	start_rev, 
    	start_RC,
	cnt_up,

	ready_par, 
	ready_rot, 
	ready_per, 
	ready_rev, 
	ready_RC,
	co
);

  input clk, rst, start_par, start_rot, start_per, start_rev, start_RC, cnt_up;
  output ready_par, ready_rot, ready_per, ready_rev, ready_RC, co;
  wire [0:4]loop_num;


  col_parity cpar(clk, rst, start_par, ready_par);

  rotate rott(clk, rst, start_rot, ready_rot);

  permute perm(clk, rst, start_per, ready_per);

  revaluate reval(clk, rst, start_rev, ready_rev);

  addRC addrc(clk, rst, start_RC, loop_num, ready_RC);

  counter24 cntr(clk, rst, cnt_up, co, loop_num);
  
 
  
endmodule

