
module dcder(
    i,
    shift_out
);
    input[0:4] i;
    output reg[0:5] shift_out;
    //output reg[0:4] to25_out;

    assign shift_out = (i == 5'd0) ? 6'd21:
		(i == 5'd1 ) ? 6'd8:
		(i == 5'd2 ) ? 6'd41:
		(i == 5'd3 ) ? 6'd45:
		(i == 5'd4 ) ? 6'd15:
		(i == 5'd5 ) ? 6'd56:
		(i == 5'd6 ) ? 6'd14:
		(i == 5'd7 ) ? 6'd18:
		(i == 5'd8 ) ? 6'd2:
		(i == 5'd9 ) ? 6'd61:
		(i == 5'd10 ) ? 6'd28:
		(i == 5'd11) ? 6'd27:
		(i == 5'd12) ? 6'd0:
		(i == 5'd13) ? 6'd1:
		(i == 5'd14) ? 6'd62:
		(i == 5'd15) ? 6'd55:
		(i == 5'd16) ? 6'd20:
		(i == 5'd17) ? 6'd36:
		(i == 5'd18) ? 6'd44:
		(i == 5'd19) ? 6'd6:
		(i == 5'd20) ? 6'd25:
		(i == 5'd21) ? 6'd39:
		(i == 5'd22) ? 6'd3:
		(i == 5'd23) ? 6'd10:
		(i == 5'd24) ? 6'd43: 6'd0;

    /*assign to25_out = (i == 3'd3 && j == 3'd3) ? 5'd0:
		(i == 3'd4 && j == 3'd3) ? 5'd1:
		(i == 3'd0 && j == 3'd3) ? 5'd2:
		(i == 3'd1 && j == 3'd3) ? 5'd3:
		(i == 3'd2 && j == 3'd3) ? 5'd4:
		(i == 3'd3 && j == 3'd4) ? 5'd5:
		(i == 3'd4 && j == 3'd4) ? 5'd6:
		(i == 3'd0 && j == 3'd4) ? 5'd7:
		(i == 3'd1 && j == 3'd4) ? 5'd8:
		(i == 3'd2 && j == 3'd4) ? 5'd9:
		(i == 3'd3 && j == 3'd0) ? 5'd10:
		(i == 3'd4 && j == 3'd0) ? 5'd11:
		(i == 3'd0 && j == 3'd0) ? 5'd12:
		(i == 3'd1 && j == 3'd0) ? 5'd13:
		(i == 3'd2 && j == 3'd0) ? 5'd14:
		(i == 3'd3 && j == 3'd1) ? 5'd15:
		(i == 3'd4 && j == 3'd1) ? 5'd16:
		(i == 3'd0 && j == 3'd1) ? 5'd17:
		(i == 3'd1 && j == 3'd1) ? 5'd18:
		(i == 3'd2 && j == 3'd1) ? 5'd19:
		(i == 3'd3 && j == 3'd2) ? 5'd20:
		(i == 3'd4 && j == 3'd2) ? 5'd21:
		(i == 3'd0 && j == 3'd2) ? 5'd22:
		(i == 3'd1 && j == 3'd2) ? 5'd23:
		(i == 3'd2 && j == 3'd2) ? 5'd24: 5'd0;
		*/
    
endmodule
    

 